----library ieee;--
--use ieee.std_logic1164.all;
--use IEEE.NUMERIC_STD.ALL;
--use STD.textio.all;
--use ieee.std_logic_textio.all;
--
--
---- Declare the Component under test
--
--entity g04_MAC_tb is
--port ( x			: in std_logic_vector(7 downto 0); -- first input
--		 y			: in std_logic_vector(8 downto 0); -- second input
--		 N			: in std_logic_vector(9 downto 0); -- total number of inputs
--		 clk		: in std_logic; --clock
--		 rst 		: in std_logic; --asynchronous active - high reset
--		 mac		: out std_logic_vector(16 downto 0); -- output of MAC unit
--		 ready 	: out std_logic); -- denotes the validity of the mac signal
--end g04_MAC_tb;
--
---- Testbench internal signals
--file file_VECTORS_X : text;
--file file_VECTORS_X : text;
--file file_RESULTS : text;
--
--constant clk_peiod : time := 100 ns;
--
--signal x_in		: in std_logic_vector(?? downto 0); 
--signal y_in			: in std_logic_vector(?? downto 0); 
--signal N_in		: in std_logic_vector(9 downto 0); 
--signal clk_in		: in std_logic; 
--signal rst_in 		: in std_logic; 
--signal mac_in		: out std_logic_vector(?? downto 0); 
--signal ready_in 	: out std_logic);
--
--
--architecture test of g04_MAC_b is
--
--begin
--
---- instantiate MAC
--	g04_MAC_INST : g04_MAC;
--	port map (x => x_in;
--				 y => y_in;
--				 N => N_in;
--				 clk => clk_in;
--				 rst => rst_in;
--				 mac => mac_out;
--				 readyS => read_out);


--	clk_generation